module Graphic_controller(input logic A,input logic B, output logic C);
assign C = A|B;
endmodule